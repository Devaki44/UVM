interface intf;
  
  bit a;
  bit b;
  bit out;
  
endinterface
