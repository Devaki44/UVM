interface intf;
  
  logic a;
  logic b;
  logic out;
  
endinterface
