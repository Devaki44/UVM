interface interf;
  bit a,b,cin;
  bit sum,cout;
endinterface
