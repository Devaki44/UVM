interface interf;
  bit clk;
  bit rst;
  bit d;
  bit q;
endinterface

